library ieee;
use ieee.std_logic_1164.all;

entity microcode is
	port (
		Address : in std_logic_vector(8 downto 0);
		Data : out std_logic_vector(23 downto 0)
	);
end microcode;

architecture impl of microcode is
begin
    PROCESS(all)
      BEGIN
         CASE (Address) IS
            WHEN "000000000" => Data <= "100000000000000000000000";
            WHEN "000001010" => Data <= "101001100000000101100100";
            WHEN "000010010" => Data <= "001000100000010001100100";
            WHEN "000010100" => Data <= "001000100000010101100100";
            WHEN "000010101" => Data <= "000000000000000000000011";
            WHEN "000010110" => Data <= "100001100000000101100111";
            WHEN "000011001" => Data <= "000000000000000000000010";
            WHEN "000011010" => Data <= "100001100000000101100110";
            WHEN "000100010" => Data <= "001000100000010001100100";
            WHEN "000100100" => Data <= "001000100000010101100100";
            WHEN "000100101" => Data <= "100000100000011000010111";
            WHEN "000101001" => Data <= "100000100000011000010110";
            WHEN "000110010" => Data <= "001000100000001001100100";
            WHEN "000110100" => Data <= "101000100000001101100100";
            WHEN "000111010" => Data <= "001000100000010001100100";
            WHEN "000111011" => Data <= "100001100000000110010100";
            WHEN "001000010" => Data <= "001000100000010001100100";
            WHEN "001000011" => Data <= "100000100000011100010100";
            WHEN "001001000" => Data <= "100001100000000100011000";
            WHEN "001010000" => Data <= "100001100000000100011100";
            WHEN "001011000" => Data <= "000001100000001100111000";
            WHEN "001011001" => Data <= "000010000001000000110100";
            WHEN "001011010" => Data <= "100001100000001000101000";
            WHEN "001100000" => Data <= "000001100000001100111100";
            WHEN "001100001" => Data <= "000010000001100000110100";
            WHEN "001100010" => Data <= "100001100000001000101100";
            WHEN "001101010" => Data <= "001000100000010001100100";
            WHEN "001101011" => Data <= "100001100000000001000000";
            WHEN "001110000" => Data <= "100001100000000000010000";
            WHEN "001111010" => Data <= "001000100000010001100100";
            WHEN "001111011" => Data <= "100001100000100001000000";
            WHEN "010000000" => Data <= "100001100000100000010000";
            WHEN "010001010" => Data <= "001000100000010001100100";
            WHEN "010001011" => Data <= "100001100001000001000000";
            WHEN "010010000" => Data <= "100001100001000000010000";
            WHEN "010011010" => Data <= "001000100000010001100100";
            WHEN "010011011" => Data <= "100001100001100001000000";
            WHEN "010100000" => Data <= "100001100001100000010000";
            WHEN "010101010" => Data <= "001000100000010001100100";
            WHEN "010101011" => Data <= "100001100010000001000000";
            WHEN "010110000" => Data <= "100001100010000000010000";
            WHEN "010111010" => Data <= "001000100000010001100100";
            WHEN "010111011" => Data <= "100001100010100001000000";
            WHEN "011000000" => Data <= "100001100010100000010000";
            WHEN "011001010" => Data <= "001000100000010001100100";
            WHEN "011001011" => Data <= "100001100011000001000000";
            WHEN "011010000" => Data <= "100001100011000000010000";
            WHEN "011011010" => Data <= "001000100000010001100100";
            WHEN "011011011" => Data <= "100001000011100001000000";
            WHEN "011100000" => Data <= "100001000011100000010000";
            WHEN "011101010" => Data <= "001000100000010001100100";
            WHEN "011101100" => Data <= "001000100000010101100100";
            WHEN "011101101" => Data <= "110000000000100000000000";
            WHEN "011110000" => Data <= "110000000000000000000000";
            WHEN "011111010" => Data <= "010000000001000001100100";
            WHEN "011111011" => Data <= "101000000000000000000000";
            WHEN "100000010" => Data <= "001000100000010001100100";
            WHEN "100000011" => Data <= "000010000000100000000000";
            WHEN "100000100" => Data <= "110000000001000001000100";
            WHEN "100001010" => Data <= "001000100000010001100100";
            WHEN "100001011" => Data <= "000010000000000000000000";
            WHEN "100001100" => Data <= "110000000001000001000100";
            WHEN "100010001" => Data <= "000000100000010000000100";
            WHEN "100010010" => Data <= "100001100000000110010100";
            WHEN "100011001" => Data <= "000000100000010000000100";
            WHEN "100011010" => Data <= "100000100000011100010100";
            WHEN "100100000" => Data <= "000000001000000000000000";
            WHEN "100100001" => Data <= "100000100000011000010101";
            WHEN "100101001" => Data <= "000000000000000000000001";
            WHEN "100101010" => Data <= "100000111000000101100101";
            WHEN "100110010" => Data <= "001000100000010001100100";
            WHEN "100110100" => Data <= "001000101000010101100100";
            WHEN "100110101" => Data <= "000000101000011001110101";
            WHEN "100110110" => Data <= "000000100000011010000101";
            WHEN "100110111" => Data <= "110000000000100000000000";
            WHEN "100111001" => Data <= "000000000000000000000001";
            WHEN "100111010" => Data <= "000000111000010001100101";
            WHEN "100111011" => Data <= "000000000000000000000001";
            WHEN "100111100" => Data <= "000000111000010101100101";
            WHEN "100111101" => Data <= "110000000000100000000000";
            WHEN "101000001" => Data <= "000100000000000000000000";
            WHEN "101001000" => Data <= "100001100100000000010000";
            WHEN "101010000" => Data <= "100001100100100000010000";
            WHEN "101011000" => Data <= "100001100101000000010000";
            WHEN OTHERS => Data <= (OTHERS => '0');
         END CASE;
      END PROCESS;
end impl;
